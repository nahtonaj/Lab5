module sext();

endmodule