module pc(RESET, PC, NEXT_PC);


endmodule