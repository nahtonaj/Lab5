module muxPC(H, MP, NextPC, ADD, HALT, PC);
endmodule